library verilog;
use verilog.vl_types.all;
entity mips_cpu is
    port(
        CLOCK_50        : in     vl_logic;
        KEY             : in     vl_logic_vector(3 downto 0);
        SW              : in     vl_logic_vector(17 downto 0);
        HEX7            : out    vl_logic_vector(6 downto 0);
        HEX6            : out    vl_logic_vector(6 downto 0);
        HEX5            : out    vl_logic_vector(6 downto 0);
        HEX4            : out    vl_logic_vector(6 downto 0);
        HEX3            : out    vl_logic_vector(6 downto 0);
        HEX2            : out    vl_logic_vector(6 downto 0);
        HEX1            : out    vl_logic_vector(6 downto 0);
        HEX0            : out    vl_logic_vector(6 downto 0);
        LEDG            : out    vl_logic_vector(7 downto 0);
        LEDR            : out    vl_logic_vector(17 downto 0);
        DRAM_ADDR       : out    vl_logic_vector(11 downto 0);
        DRAM_BA_0       : out    vl_logic;
        DRAM_BA_1       : out    vl_logic;
        DRAM_CAS_N      : out    vl_logic;
        DRAM_CKE        : out    vl_logic;
        DRAM_CLK        : out    vl_logic;
        DRAM_CS_N       : out    vl_logic;
        DRAM_DQ         : inout  vl_logic_vector(15 downto 0);
        DRAM_LDQM       : out    vl_logic;
        DRAM_UDQM       : out    vl_logic;
        DRAM_RAS_N      : out    vl_logic;
        DRAM_WE_N       : out    vl_logic;
        FL_ADDR         : out    vl_logic_vector(21 downto 0);
        FL_DQ           : inout  vl_logic_vector(7 downto 0);
        FL_CE_N         : out    vl_logic;
        FL_OE_N         : out    vl_logic;
        FL_RST_N        : out    vl_logic;
        FL_WE_N         : out    vl_logic;
        SRAM_ADDR       : out    vl_logic_vector(17 downto 0);
        SRAM_DQ         : inout  vl_logic_vector(15 downto 0);
        SRAM_UB_N       : out    vl_logic;
        SRAM_LB_N       : out    vl_logic;
        SRAM_WE_N       : out    vl_logic;
        SRAM_OE_N       : out    vl_logic;
        SRAM_CE_N       : out    vl_logic
    );
end mips_cpu;
