library verilog;
use verilog.vl_types.all;
entity test_bp is
end test_bp;
