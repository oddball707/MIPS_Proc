library verilog;
use verilog.vl_types.all;
entity iq is
end iq;
