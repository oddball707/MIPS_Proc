library verilog;
use verilog.vl_types.all;
entity test_mips_cpu is
end test_mips_cpu;
